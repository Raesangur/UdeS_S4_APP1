14 gid=414328
14 uid=414328
27 mtime=1651691362.486951
