s <=  a xor b  xor c;
r <= (a and b) or (a and c) or (c and b);
