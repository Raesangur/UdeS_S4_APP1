14 gid=414328
14 uid=414328
26 mtime=1651691361.91994
